* Simple Resistive Attenuator (Voltage Divider)

Vin IN 0 SIN(0 10 1k)

R1 IN OUT 10k
R2 OUT 0 10k

.control
set filetype=ascii
tran 0.1ms 5ms
write attenuator.raw
.endc

.end
