* Half Wave Rectifier

Vin IN 0 SIN(0 10 1k)

D1 IN OUT Dmodel
Rload OUT 0 1k

.model Dmodel D(Is=1e-14 N=1)

.control
set filetype=ascii
tran 0.1ms 5ms
write rectifier.raw
.endc

.end
