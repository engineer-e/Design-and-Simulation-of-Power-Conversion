* Title : Simple attenuator circuit

* Netlist
V1 a 0 100v
R1 a b 20
R2 b 0 10

* Control commands
.control
op
print v(a) v(b) v(a,b) i(v1)
.endc
.end