* Title : Half wave rectifier

* Netlist

V1 a 0 sin(0 100 50 0 0)
D1 a c dmodel
R1 c b 10
R2 b 0 10

* Model 
.model dmodel D()

* Control
.control 
set color0 = white ; set background color white
set color1 = black ; set foreground color black
tran 1us 40ms uic
plot v(a) v(b)
.endc
.end