* Half Wave Rectifier

Vin IN 0 SIN(0 100 50 0 0)

D1 IN OUT Dmodel
Rload OUT 0 1k

.model Dmodel D(Is=1e-14 N=1)

.control
set filetype=ascii
tran 0.1ms 40ms
write half-wave-rectifier.raw
.endc

.end
